/*
 
 
 
 */

module ExecuteTwo
  (
   input logic clk,
   input logic rstn
   );


endmodule // ExecuteTwo
