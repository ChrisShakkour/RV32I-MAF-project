/*
 
 
 
 */

module IDMemory
  (
   input logic clk,
   input logic rstn
   );


endmodule // IDMemory
