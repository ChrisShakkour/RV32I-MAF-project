// all the OP_CODE of Flot instructions 
