/*
 
 
 
 */

module LoadStore 
  (
   input logic         clk,
   input logic         rstn,
   
);

endmodule
