/*
 
 
 
 
 */

module InstructionFetch 
  (
   input logic clk,
   input logic rstn
   );





endmodule // InstructionFetch
