/*
 
 
 
 */

module WriteBack
  (
   input logic clk,
   input logic rstn
   );



endmodule // WriteBack
