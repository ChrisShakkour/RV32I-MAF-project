/*
 
 
 
 */

module Decode
  (
   input logic clk,
   input logic rstn
   );



endmodule // Decode
