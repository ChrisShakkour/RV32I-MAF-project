/*
 
 
 
 */

module ExecuteOne 
  (
   input logic clk,
   input logic rstn
   );


endmodule // ExecuteOne

   
